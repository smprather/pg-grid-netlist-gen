.subckt BUFX12 A Y VDD VSS
.ends
