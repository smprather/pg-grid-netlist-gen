.subckt DCAPX32 VDD VSS
.ends
